module(
    input logic clk,
    input logic n_rst,
    input logic hsel,
    input logic [3:0] haddr,
    input logic hsize,
    input logic htrans[1:0],
    input logic hwrite,
    input logic hwdata[15:0],
    output logic hrdata[15:0],
    output logic hresp
);



endmodule